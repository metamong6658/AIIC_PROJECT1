`timescale 1ns/1ns
`include "Controller.v"
`include "PE.v"
`include "RAM.v"
`include "ReLu.v"
`include "Sigmoid.v"
`include "ROM.v"

module tb_Controller;
parameter Qw = 122;
parameter sigmoid_max = 1874;
parameter TESTNUMBER = 20;
parameter ROM0_ADDR_MAX = 67280;
parameter ROM0_ADDR_WIDTH = 17;
parameter INFILE0 = "RTL_test_data.hex";
parameter INFILE1 = "weights_layer1.hex";
parameter INFILE2 = "weights_layer2.hex";
parameter INFILE3 = "weights_layer3.hex";
parameter INFILE4 = "weights_layer4.hex";
localparam [19:0] LABEL =           20'b10011_00110_00000_11000;
localparam [19:0] SWPREDICTION =    20'b10011_00110_00000_11000; // 100%
reg i_clk;
reg i_rst;
reg i_en;
wire [19:0] o_array; // 60%
wire done;

Controller #(
    .Qw(Qw), 
    .sigmoid_max(sigmoid_max),
    .TESTNUMBER(TESTNUMBER),
    .ROM0_ADDR_MAX(ROM0_ADDR_MAX),
    .ROM0_ADDR_WIDTH(ROM0_ADDR_WIDTH),
    .INFILE0(INFILE0),
    .INFILE1(INFILE1),
    .INFILE2(INFILE2),
    .INFILE3(INFILE3),
    .INFILE4(INFILE4)
    ) i_Controller(
    .i_clk(i_clk),
    .i_rst(i_rst),
    .i_en(i_en),
    .o_array(o_array),
    .done(done)
);

always #5 i_clk = ~i_clk;

initial begin
    i_clk = 0;
    i_rst = 0;
    i_en = 0;
    #10;
    i_rst = 1;
    #10;
    i_rst = 0;
    #10;
    i_en = 1;
    // TEST1
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST2
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST3
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST4
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST5
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST6
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST7
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST8
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST9
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST10
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST1
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST2
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST3
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST4
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST5
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST6
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST7
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST8
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST9
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    // TEST10
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    #1000000;
    $finish;
end

endmodule